******
*==
v1 1 0 2
v2 2 0 3
r1 1 2 1
.dc v1 1 2 0.5
.end
